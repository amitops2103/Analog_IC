** sch_path: /home/amitvlsi01/untitled-1.sch
.subckt untitled-1 VDD A Y GND
*.PININFO A:I VDD:I GND:I Y:O
XM1 Y A GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
**** begin user architecture code
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
**** end user architecture code
.ends
