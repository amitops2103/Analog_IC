.TITLE Diode Experiment

*.MODEL dio1 D (bv=50 is=1e-13 n=1.05)


D1    vin    vout   dio1
R1    vout   GND    1k
*C1    vout   GND    1p

Vs    vin   GND    0 SIN(0 1 1e3 0 0 0 )
.MODEL dio1 D (bv=50 is=1e-13 n=1.05)
.OP
.TRAN 1u 4m

.END

